`define HEADER 8
`define PARITY 8
`define payload 8